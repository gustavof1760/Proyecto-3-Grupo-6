`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    19:00:46 05/10/2017
// Design Name: 
// Module Name:    Temporizador 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Temporizador(clk, reset, carga_temp, temp_sel, listo);

/////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
////ENTRADAS y SALIDAS
/////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
input clk, reset, carga_temp;
input [1:0] temp_sel;
output listo;

/////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
//// Registros
/////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////	

reg [3:0] contador;
reg [3:0] contador_sig;
reg listo;

/////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
/////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////	
parameter [3:0] Ts_ad = 4'd3;
parameter [3:0] Tc_ac = 4'd7;
parameter [3:0] Tw = 4'd12;
/////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
/////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
//Registro de estado

//Logica de contador Siguiente
always@(reset or carga_temp or temp_sel or listo or contador) 
    begin
        casex({reset, carga_temp, temp_sel, listo})
        5'b1xxxx: contador_sig = 4'b0;
        5'b0101x: contador_sig = Ts_ad;
        5'b0110x: contador_sig = Tc_ac;
        5'b0111x: contador_sig = Tw;
        5'b00xx0: contador_sig = contador - 1'b1;
        5'b00xx1: contador_sig = contador;
        default: contador_sig = contador;
        endcase
    end

always @(posedge clk) 
    begin
         contador <= contador_sig;
    end

always @* 
    begin
        listo = !(|contador) ; //Cuenta terminada
    end
	
endmodule